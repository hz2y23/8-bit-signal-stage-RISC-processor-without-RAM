
`define ADD 	3'b000
`define SLLI  	3'b001
`define J	 	3'b010
`define SUB 	3'b011
`define BLT		3'b100
`define ADDI 	3'b101
`define SRL 	3'b110
`define BEQ		3'b111