
`define RADD 		3'b000
`define RSLL 		3'b001
`define RSUB		3'b010
`define RSRL 		3'b011
`define NOP 		3'b100